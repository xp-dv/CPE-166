/* Traffic Signal Color Package */
package traffic_signal_colors_pkg;
  // 0 = Flashing Red
  // 1 = Red
  // 2 = Yellow
  // 3 = Green
  typedef enum logic [1:0] {FLASHING, RED, YELLOW, GREEN} color_e;
endpackage

