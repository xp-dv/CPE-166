/* Datapath Top-Level Module */
module datapath(
  input clr, clk, cin;
  input [3:0] m0, m1, m2;
  input [2:0] w;
  input [3:0] ce;
  input [1:0] sel;
  input [2:0] s;
  output [3:0] r0, r1, r2;
);



endmodule
