---- Watch Block ----
