---- Stopwatch Test Bench ----
